module CosTable(
  input  [7:0] cos_ad, // 読み込みアドレス
  output signed [7:0] cos_rd  // 読み込みデータ
);
  reg signed [7:0] cos[256]={
     64, 64, 64, 64, 64, 64, 63, 63, 63, 62, 62, 62, 61, 61, 60, 60,
     59, 59, 58, 57, 56, 56, 55, 54, 53, 52, 51, 50, 49, 48, 47, 46,
     45, 44, 43, 42, 41, 39, 38, 37, 36, 34, 33, 32, 30, 29, 27, 26,
     24, 23, 22, 20, 19, 17, 16, 14, 12, 11,  9,  8,  6,  5,  3,  2,
      0, -2, -3, -5, -6, -8, -9,-11,-12,-14,-16,-17,-19,-20,-22,-23,
    -24,-26,-27,-29,-30,-32,-33,-34,-36,-37,-38,-39,-41,-42,-43,-44,
    -45,-46,-47,-48,-49,-50,-51,-52,-53,-54,-55,-56,-56,-57,-58,-59,
    -59,-60,-60,-61,-61,-62,-62,-62,-63,-63,-63,-64,-64,-64,-64,-64,
    -64,-64,-64,-64,-64,-64,-63,-63,-63,-62,-62,-62,-61,-61,-60,-60,
    -59,-59,-58,-57,-56,-56,-55,-54,-53,-52,-51,-50,-49,-48,-47,-46,
    -45,-44,-43,-42,-41,-39,-38,-37,-36,-34,-33,-32,-30,-29,-27,-26,
    -24,-23,-22,-20,-19,-17,-16,-14,-12,-11, -9, -8, -6, -5, -3, -2,
      0,  2,  3,  5,  6,  8,  9, 11, 12, 14, 16, 17, 19, 20, 22, 23,
     24, 26, 27, 29, 30, 32, 33, 34, 36, 37, 38, 39, 41, 42, 43, 44,
     45, 46, 47, 48, 49, 50, 51, 52, 53, 54, 55, 56, 56, 57, 58, 59,
     59, 60, 60, 61, 61, 62, 62, 62, 63, 63, 63, 64, 64, 64, 64, 64
  }; // ラインバッファ 256ドット*2ライン
  assign cos_rd = cos[cos_ad]; // 読み込み
endmodule


module StartTable(
  input  [7:0] sta_ad, // 読み込みアドレス
  output [31:0] sta_rd  // 読み込みデータ
);
  assign sta_rd = sta[sta_ad]; // 読み込み
//  reg [31:0] sta2[1:0]='{32'h00000800,{16'hff40,16'h0400}};

  reg [31:0] sta[256]={
    32'h00000800,{16'hff40,16'h0900},{16'hfee0,16'h0980},{16'hfe20,16'h0a80},{16'hfdc0,16'h0b00},{16'hfd00,16'h0c00},{16'hfd20,16'h0ce0},{16'hfc60,16'h0de0},{16'hfc00,16'h0e60},{16'hfbc0,16'h0fc0},{16'hfb00,16'h10c0},{16'hfaa0,16'h1140},{16'hfa60,16'h12a0},{16'hfa00,16'h1320},{16'hf9c0,16'h1480},{16'hf960,16'h1500},
    {16'hf980,16'h15e0},{16'hf8c0,16'h16e0},{16'hf8e0,16'h17c0},{16'hf8a0,16'h1920},{16'hf8c0,16'h1a00},{16'hf800,16'h1b00},{16'hf820,16'h1be0},{16'hf840,16'h1cc0},{16'hf800,16'h1e20},{16'hf820,16'h1f00},{16'hf840,16'h1fe0},{16'hf860,16'h20c0},{16'hf820,16'h2220},{16'hf840,16'h2300},{16'hf860,16'h23e0},{16'hf880,16'h24c0},
    {16'hf8a0,16'h25a0},{16'hf8c0,16'h2680},{16'hf8e0,16'h2760},{16'hf900,16'h2840},{16'hf920,16'h2920},{16'hf9c0,16'h2a60},{16'hf9e0,16'h2b40},{16'hfa00,16'h2c20},{16'hfa20,16'h2d00},{16'hfac0,16'h2e40},{16'hfae0,16'h2f20},{16'hfb00,16'h3000},{16'hfc00,16'h30c0},{16'hfc20,16'h31a0},{16'hfcc0,16'h32e0},{16'hfce0,16'h33c0},
    {16'hfde0,16'h3480},{16'hfe00,16'h3560},{16'hfe80,16'h35c0},{16'hff20,16'h3700},{16'hffa0,16'h3760},{16'h0040,16'h38a0},{16'h00c0,16'h3900},{16'h01c0,16'h39c0},{16'h0260,16'h3b00},{16'h02e0,16'h3b60},{16'h03e0,16'h3c20},{16'h0400,16'h3d00},{16'h0500,16'h3dc0},{16'h0580,16'h3e20},{16'h0680,16'h3ee0},{16'h0700,16'h3f40},
    {16'h0800,16'h4000},{16'h0900,16'h40c0},{16'h0980,16'h4120},{16'h0a80,16'h41e0},{16'h0b00,16'h4240},{16'h0c00,16'h4300},{16'h0ce0,16'h42e0},{16'h0de0,16'h43a0},{16'h0e60,16'h4400},{16'h0fc0,16'h4440},{16'h10c0,16'h4500},{16'h1140,16'h4560},{16'h12a0,16'h45a0},{16'h1320,16'h4600},{16'h1480,16'h4640},{16'h1500,16'h46a0},
    {16'h15e0,16'h4680},{16'h16e0,16'h4740},{16'h17c0,16'h4720},{16'h1920,16'h4760},{16'h1a00,16'h4740},{16'h1b00,16'h4800},{16'h1be0,16'h47e0},{16'h1cc0,16'h47c0},{16'h1e20,16'h4800},{16'h1f00,16'h47e0},{16'h1fe0,16'h47c0},{16'h20c0,16'h47a0},{16'h2220,16'h47e0},{16'h2300,16'h47c0},{16'h23e0,16'h47a0},{16'h24c0,16'h4780},
    {16'h25a0,16'h4760},{16'h2680,16'h4740},{16'h2760,16'h4720},{16'h2840,16'h4700},{16'h2920,16'h46e0},{16'h2a60,16'h4640},{16'h2b40,16'h4620},{16'h2c20,16'h4600},{16'h2d00,16'h45e0},{16'h2e40,16'h4540},{16'h2f20,16'h4520},{16'h3000,16'h4500},{16'h30c0,16'h4400},{16'h31a0,16'h43e0},{16'h32e0,16'h4340},{16'h33c0,16'h4320},
    {16'h3480,16'h4220},{16'h3560,16'h4200},{16'h35c0,16'h4180},{16'h3700,16'h40e0},{16'h3760,16'h4060},{16'h38a0,16'h3fc0},{16'h3900,16'h3f40},{16'h39c0,16'h3e40},{16'h3b00,16'h3da0},{16'h3b60,16'h3d20},{16'h3c20,16'h3c20},{16'h3d00,16'h3c00},{16'h3dc0,16'h3b00},{16'h3e20,16'h3a80},{16'h3ee0,16'h3980},{16'h3f40,16'h3900},
    {16'h4000,16'h3800},{16'h40c0,16'h3700},{16'h4120,16'h3680},{16'h41e0,16'h3580},{16'h4240,16'h3500},{16'h4300,16'h3400},{16'h42e0,16'h3320},{16'h43a0,16'h3220},{16'h4400,16'h31a0},{16'h4440,16'h3040},{16'h4500,16'h2f40},{16'h4560,16'h2ec0},{16'h45a0,16'h2d60},{16'h4600,16'h2ce0},{16'h4640,16'h2b80},{16'h46a0,16'h2b00},
    {16'h4680,16'h2a20},{16'h4740,16'h2920},{16'h4720,16'h2840},{16'h4760,16'h26e0},{16'h4740,16'h2600},{16'h4800,16'h2500},{16'h47e0,16'h2420},{16'h47c0,16'h2340},{16'h4800,16'h21e0},{16'h47e0,16'h2100},{16'h47c0,16'h2020},{16'h47a0,16'h1f40},{16'h47e0,16'h1de0},{16'h47c0,16'h1d00},{16'h47a0,16'h1c20},{16'h4780,16'h1b40},
    {16'h4760,16'h1a60},{16'h4740,16'h1980},{16'h4720,16'h18a0},{16'h4700,16'h17c0},{16'h46e0,16'h16e0},{16'h4640,16'h15a0},{16'h4620,16'h14c0},{16'h4600,16'h13e0},{16'h45e0,16'h1300},{16'h4540,16'h11c0},{16'h4520,16'h10e0},{16'h4500,16'h1000},{16'h4400,16'h0f40},{16'h43e0,16'h0e60},{16'h4340,16'h0d20},{16'h4320,16'h0c40},
    {16'h4220,16'h0b80},{16'h4200,16'h0aa0},{16'h4180,16'h0a40},{16'h40e0,16'h0900},{16'h4060,16'h08a0},{16'h3fc0,16'h0760},{16'h3f40,16'h0700},{16'h3e40,16'h0640},{16'h3da0,16'h0500},{16'h3d20,16'h04a0},{16'h3c20,16'h03e0},{16'h3c00,16'h0300},{16'h3b00,16'h0240},{16'h3a80,16'h01e0},{16'h3980,16'h0120},{16'h3900,16'h00c0},
    {16'h3800,16'h0000},{16'h3700,16'hff40},{16'h3680,16'hfee0},{16'h3580,16'hfe20},{16'h3500,16'hfdc0},{16'h3400,16'hfd00},{16'h3320,16'hfd20},{16'h3220,16'hfc60},{16'h31a0,16'hfc00},{16'h3040,16'hfbc0},{16'h2f40,16'hfb00},{16'h2ec0,16'hfaa0},{16'h2d60,16'hfa60},{16'h2ce0,16'hfa00},{16'h2b80,16'hf9c0},{16'h2b00,16'hf960},
    {16'h2a20,16'hf980},{16'h2920,16'hf8c0},{16'h2840,16'hf8e0},{16'h26e0,16'hf8a0},{16'h2600,16'hf8c0},{16'h2500,16'hf800},{16'h2420,16'hf820},{16'h2340,16'hf840},{16'h21e0,16'hf800},{16'h2100,16'hf820},{16'h2020,16'hf840},{16'h1f40,16'hf860},{16'h1de0,16'hf820},{16'h1d00,16'hf840},{16'h1c20,16'hf860},{16'h1b40,16'hf880},
    {16'h1a60,16'hf8a0},{16'h1980,16'hf8c0},{16'h18a0,16'hf8e0},{16'h17c0,16'hf900},{16'h16e0,16'hf920},{16'h15a0,16'hf9c0},{16'h14c0,16'hf9e0},{16'h13e0,16'hfa00},{16'h1300,16'hfa20},{16'h11c0,16'hfac0},{16'h10e0,16'hfae0},{16'h1000,16'hfb00},{16'h0f40,16'hfc00},{16'h0e60,16'hfc20},{16'h0d20,16'hfcc0},{16'h0c40,16'hfce0},
    {16'h0b80,16'hfde0},{16'h0aa0,16'hfe00},{16'h0a40,16'hfe80},{16'h0900,16'hff20},{16'h08a0,16'hffa0},{16'h0760,16'h0040},{16'h0700,16'h00c0},{16'h0640,16'h01c0},{16'h0500,16'h0260},{16'h04a0,16'h02e0},{16'h03e0,16'h03e0},{16'h0300,16'h0400},{16'h0240,16'h0500},{16'h01e0,16'h0580},{16'h0120,16'h0680},{16'h00c0,16'h0700}
  };
endmodule
